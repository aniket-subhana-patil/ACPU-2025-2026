library IEEE;
use IEEE.std_logic_1164.ALL;
use IEEE.numeric_std.ALL;

-- TODO include your package

entity memory is
	generic (
		-- TODO declare generics word_size and mem_size
	);
	port (
		-- TODO declare ports addr_write, addr_read, data_write, data_read, writen_en, read_en, clk
	);
end entity memory;

architecture behav of memory is

	-- TODO declare types and signals

begin
 
	-- TODO add implementation

end behav;


